module TRV32I_core (
    input           clk, rst;
    input   [31:0]  inst;
    output  [31:0]  pc;
    output  [31:0]  mem_addr;
    output          mem_read_en, mem_write_en;
    output  [3:0]   write_byte_en;
    inout   [31:0]  mem_data;
);

    //datapath

    //ctlpath


endmodule
