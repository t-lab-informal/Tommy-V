module TRV32I_top #(
    parameter B_WIDTH = 32;
) (
    input           clk, rst;
    output  [31:0]  pc, inst;
    output          mem_read_en, mem_write_en;
    output  [B_WIDTH-1:0] mem_data;
);

    //datapath

    //ctlpath


endmodule
